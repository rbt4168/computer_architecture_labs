module AndUnit (
    input value_a, value_b,
    output value_o
);
    assign value_o = value_a & value_b;
endmodule